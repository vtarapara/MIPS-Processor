module and_32_bitwise(a, b, res);
    input [31:0] a;
    input [31:0] b;
    output [31:0] res;

    and and_gate0(res[0], a[0], b[0]);
    and and_gate1(res[1], a[1], b[1]);
    and and_gate2(res[2], a[2], b[2]);
    and and_gate3(res[3], a[3], b[3]);
    and and_gate4(res[4], a[4], b[4]);
    and and_gate5(res[5], a[5], b[5]);
    and and_gate6(res[6], a[6], b[6]);
    and and_gate7(res[7], a[7], b[7]);
    and and_gate8(res[8], a[8], b[8]);
    and and_gate9(res[9], a[9], b[9]);
    and and_gate10(res[10], a[10], b[10]);
    and and_gate11(res[11], a[11], b[11]);
    and and_gate12(res[12], a[12], b[12]);
    and and_gate13(res[13], a[13], b[13]);
    and and_gate14(res[14], a[14], b[14]);
    and and_gate15(res[15], a[15], b[15]);
    and and_gate16(res[16], a[16], b[16]);
    and and_gate17(res[17], a[17], b[17]);
    and and_gate18(res[18], a[18], b[18]);
    and and_gate19(res[19], a[19], b[19]);
    and and_gate20(res[20], a[20], b[20]);
    and and_gate21(res[21], a[21], b[21]);
    and and_gate22(res[22], a[22], b[22]);
    and and_gate23(res[23], a[23], b[23]);
    and and_gate24(res[24], a[24], b[24]);
    and and_gate25(res[25], a[25], b[25]);
    and and_gate26(res[26], a[26], b[26]);
    and and_gate27(res[27], a[27], b[27]);
    and and_gate28(res[28], a[28], b[28]);
    and and_gate29(res[29], a[29], b[29]);
    and and_gate30(res[30], a[30], b[30]);
    and and_gate31(res[31], a[31], b[31]);
    
endmodule

