module not_32_bitwise(a, res);
    input [31:0] a;
    output [31:0] res;

    not not_gate0(res[0], a[0]);
    not not_gate1(res[1], a[1]);
    not not_gate2(res[2], a[2]);
    not not_gate3(res[3], a[3]);
    not not_gate4(res[4], a[4]);
    not not_gate5(res[5], a[5]);
    not not_gate6(res[6], a[6]);
    not not_gate7(res[7], a[7]);
    not not_gate8(res[8], a[8]);
    not not_gate9(res[9], a[9]);
    not not_gate10(res[10], a[10]);
    not not_gate11(res[11], a[11]);
    not not_gate12(res[12], a[12]);
    not not_gate13(res[13], a[13]);
    not not_gate14(res[14], a[14]);
    not not_gate15(res[15], a[15]);
    not not_gate16(res[16], a[16]);
    not not_gate17(res[17], a[17]);
    not not_gate18(res[18], a[18]);
    not not_gate19(res[19], a[19]);
    not not_gate20(res[20], a[20]);
    not not_gate21(res[21], a[21]);
    not not_gate22(res[22], a[22]);
    not not_gate23(res[23], a[23]);
    not not_gate24(res[24], a[24]);
    not not_gate25(res[25], a[25]);
    not not_gate26(res[26], a[26]);
    not not_gate27(res[27], a[27]);
    not not_gate28(res[28], a[28]);
    not not_gate29(res[29], a[29]);
    not not_gate30(res[30], a[30]);
    not not_gate31(res[31], a[31]);
    
endmodule
