module register65(q, d, clk, en, clr);
    output [64:0] q;
    input [64:0] d;
    input clk;
    input en;
    input clr;
    
    // 65 bit
    dffe_ref flip_flop0(.q(q[0]), .d(d[0]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop1(.q(q[1]), .d(d[1]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop2(.q(q[2]), .d(d[2]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop3(.q(q[3]), .d(d[3]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop4(.q(q[4]), .d(d[4]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop5(.q(q[5]), .d(d[5]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop6(.q(q[6]), .d(d[6]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop7(.q(q[7]), .d(d[7]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop8(.q(q[8]), .d(d[8]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop9(.q(q[9]), .d(d[9]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop10(.q(q[10]), .d(d[10]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop11(.q(q[11]), .d(d[11]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop12(.q(q[12]), .d(d[12]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop13(.q(q[13]), .d(d[13]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop14(.q(q[14]), .d(d[14]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop15(.q(q[15]), .d(d[15]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop16(.q(q[16]), .d(d[16]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop17(.q(q[17]), .d(d[17]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop18(.q(q[18]), .d(d[18]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop19(.q(q[19]), .d(d[19]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop20(.q(q[20]), .d(d[20]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop21(.q(q[21]), .d(d[21]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop22(.q(q[22]), .d(d[22]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop23(.q(q[23]), .d(d[23]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop24(.q(q[24]), .d(d[24]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop25(.q(q[25]), .d(d[25]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop26(.q(q[26]), .d(d[26]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop27(.q(q[27]), .d(d[27]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop28(.q(q[28]), .d(d[28]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop29(.q(q[29]), .d(d[29]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop30(.q(q[30]), .d(d[30]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop31(.q(q[31]), .d(d[31]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop32(.q(q[32]), .d(d[32]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop33(.q(q[33]), .d(d[33]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop34(.q(q[34]), .d(d[34]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop35(.q(q[35]), .d(d[35]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop36(.q(q[36]), .d(d[36]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop37(.q(q[37]), .d(d[37]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop38(.q(q[38]), .d(d[38]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop39(.q(q[39]), .d(d[39]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop40(.q(q[40]), .d(d[40]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop41(.q(q[41]), .d(d[41]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop42(.q(q[42]), .d(d[42]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop43(.q(q[43]), .d(d[43]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop44(.q(q[44]), .d(d[44]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop45(.q(q[45]), .d(d[45]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop46(.q(q[46]), .d(d[46]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop47(.q(q[47]), .d(d[47]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop48(.q(q[48]), .d(d[48]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop49(.q(q[49]), .d(d[49]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop50(.q(q[50]), .d(d[50]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop51(.q(q[51]), .d(d[51]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop52(.q(q[52]), .d(d[52]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop53(.q(q[53]), .d(d[53]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop54(.q(q[54]), .d(d[54]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop55(.q(q[55]), .d(d[55]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop56(.q(q[56]), .d(d[56]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop57(.q(q[57]), .d(d[57]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop58(.q(q[58]), .d(d[58]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop59(.q(q[59]), .d(d[59]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop60(.q(q[60]), .d(d[60]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop61(.q(q[61]), .d(d[61]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop62(.q(q[62]), .d(d[62]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop63(.q(q[63]), .d(d[63]), .clk(clk), .en(en), .clr(clr));
    dffe_ref flip_flop64(.q(q[64]), .d(d[64]), .clk(clk), .en(en), .clr(clr));
endmodule